/*

Disenador: Paulina Vianney Núñez Luna
Modulo: agent_port1_pkg
Compania: Cinvestav
Contacto: paulinav.nunezl@gmail.com

*/
package agent_port1_pkg;
	import uvm_pkg::*;
	`include "uvm_macros.svh"
	
	`include "port1_monitor.svh"
	`include "port1_driver.svh"
	`include "port1_scb.svh"
	`include "port1_sqr.svh"
	`include "port1_subs.svh"
	`include "agent_port1.svh"
	
endpackage
