package ram_env_pkg;
	import uvm_pkg::*;
	`include "uvm_macros.svh"
	
	`include "ram_env.svh"
	`include "ram_scb.svh"
	
endpackage
