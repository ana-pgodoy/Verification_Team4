package ram_test_pkg;
	import uvm_pkg::*;
	import ram_env_pkg::*;	
	`include "uvm_macros.svh"
	
	`include "ram_base_test.svh"	
endpackage
