package ram_env_pkg;
	import uvm_pkg::*;
	`include "uvm_macros.svh"
	
	`include "agent_port1_pkg.sv"
	`include "agent_port0_pkg.sv"
	`include "ram_env.svh"
	`include "ram_scb.svh"
	
endpackage
