package ram_env_pkg;
	import uvm_pkg::*;
	
	import agent_port0_pkg::*;
	import agent_port1_pkg::*;
	`include "uvm_macros.svh"
	`include "ram_scb.svh"
	`include "ram_env.svh"
	
endpackage
