/*
Atribute: port0_subs
Author: Ana Paula Godoy Monroy
Date: 
Version:
File name: port0_subs.sv
*/
