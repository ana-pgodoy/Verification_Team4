class port1_read_10_seq_cs1 extends port1_base_seq;

endclass
