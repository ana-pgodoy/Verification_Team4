
class port0_read_10_seq_cs0 extends port0_base_seq;
	
endclass