/*
Atribute: port1_read_10_seq_cs1
Author: Paulina Vianney Núñez Luna
Date: 20/07/2023
Version: 1
File name: port1_read_10_seq_cs1.svh
*/

class port1_read_10_seq_cs1 extends port1_base_seq;

endclass
