/*

Disenador: Benjamin Gonzalez Alvarado
Modulo: agent_port0_pkg
Compania: Cinvestav
Contacto: a.g.ben.min@gmail.com

*/
package agent_port0_pkg;
	import uvm_pkg::*;
	`include "uvm_macros.svh"
	
	`include "port0_monitor.svh"
	`include "port0_driver.svh"
	`include "port0_scb.svh"
	`include "port0_sqr.svh"
	`include "port0_subs.svh"
	`include "agent_port0.svh"
	
endpackage
