class agent_port0 extends uvm_agent

endclass