class agent_port0 extends uvm_agent
	`uvm_component_utils(agent_port0)
endclass