package ram_defines_pkg;
  import uvm_pkg::*;
	`include "uvm_macros.svh"
//Parameters port0
  `define WMASK_WIDTH       3'h4
  `define ADDR_WIDTH        4'hA
  `define DATA_WIDTH        6'h20

//Parameters port1  
  `define ADDR_WIDTH_1      4'hA
  `define WMASK_WIDTH_1     6'h20
endpackage
