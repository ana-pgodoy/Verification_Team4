/*
Atribute: agent_port1_pkg
Author: Paulina Vianney Núñez Luna
Date: 4/07/2023
File name: agent_port1_pkg
*/
package agent_port1_pkg;
	import uvm_pkg::*;
	`include "uvm_macros.svh"
	
	`include "port1_transaction.svh"
	`include "port1_monitor.svh"
	`include "port1_driver.svh"
	`include "port1_scb.svh"
	`include "port1_seq.svh"
	`include "port1_subs.svh"
	`include "agent_port1.svh"
	
endpackage
