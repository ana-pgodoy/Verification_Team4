class agent_port0 extends uvm_agent
	`uvm_component_utils(agent_port0)
	
	
	function new(input string name, uvm_component parent);
		super.new(name,parent);
	endfunction
	
endclass